module ex

print("Hello, World!")
